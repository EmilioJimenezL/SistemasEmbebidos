module control (
    input reset,
    input clk,
    input [1:0] irq,
    output reg rw,
    input [3:0] datoin,
    output reg [7:0] pcontrol,
    input [3:0] re,
    input [7:0] pcout,
    output reg [4:0] cs
);

// Definici�n de estados - MANTENIENDO DISE�O ORIGINAL
localparam [4:0] 
    d0 = 0, d1 = 1, d2 = 2, d3 = 3, d4 = 4, d5 = 5, d6 = 6, d7 = 7, 
    d8 = 8, d9 = 9, d10 = 10, d11 = 11, d12 = 12, d13 = 13, d14 = 14, 
    d15 = 15, d16 = 16, d17 = 17;

reg [4:0] edo_presente, edo_futuro;
reg [7:0] f;

// Proceso 1: L�gica del estado futuro - COMBINACIONAL
always @(*) begin
    if (reset) begin
        edo_futuro = d0;
        pcontrol = 8'b11111111;
        rw = 1'b0;
        cs = 5'b11110;
    end else begin
        // Valores por defecto - MANTENER ESTADO ACTUAL
        edo_futuro = edo_presente;
        pcontrol = pcontrol;
        rw = rw;
        cs = cs;
        
        case (edo_presente)
            d0: begin
                if (irq == 2'b10) begin
                    cs = 5'b11100;
                    edo_futuro = d1;
                end else if (irq == 2'b01) begin
                    cs = 5'b11100;
                    edo_futuro = d1;
                end else begin
                    edo_futuro = d3;
                    cs = 5'b11111;  // ? INCREMENTAR PC - COMO EN VHDL
                end
            end
            
            d3: begin
                cs = 5'b10110;  // Leer memoria
                rw = 1'b1;
                edo_futuro = d4;
            end
            
            d4: begin
                rw = 1'b0;
                case (datoin)
                    4'b0000: begin  // CARGAR A
                        cs = 5'b00001; 
                        edo_futuro = d2;
                    end
                    4'b0001: begin  // CARGAR B
                        cs = 5'b00010; 
                        edo_futuro = d5;
                    end
                    4'b0010: begin cs = 5'b00011; edo_futuro = d5; end
                    4'b0011: begin cs = 5'b00100; edo_futuro = d5; end
                    4'b0100: begin cs = 5'b00101; edo_futuro = d5; end
                    4'b0101: begin cs = 5'b00110; edo_futuro = d5; end
                    4'b0110: begin  // STORE
                        cs = 5'b11111;  // ? INCREMENTAR PC para leer direcci�n
                        edo_futuro = d6;
                    end
                    // ... otros casos mantienen l�gica original
                    default: begin 
                        cs = 5'b11101; 
                        edo_futuro = d0; 
                    end
                endcase
            end
            
            d2: begin
                // Estado para operaciones de 1 byte
                cs = 5'b11111;  // ? INCREMENTAR PC despu�s de operaci�n
                edo_futuro = d5;
            end
            
            d5: begin
                cs = 5'b10101;
                edo_futuro = d11;
            end
            
            d6: begin
                cs = 5'b10110;  // Leer byte de direcci�n baja
                rw = 1'b1;
                edo_futuro = d12;
            end
            
            d12: begin
                cs = 5'b11111;  // ? INCREMENTAR PC para leer siguiente byte
                rw = 1'b0;
                pcontrol[3:0] = datoin;  // Guardar byte bajo
                edo_futuro = d13;
            end
            
            d13: begin
                cs = 5'b10110;  // Leer byte de direcci�n alta  
                rw = 1'b1;
                edo_futuro = d14;
            end
            
            d14: begin
                rw = 1'b0;
                cs = 5'b11010;
                pcontrol[7:4] = datoin;  // Guardar byte alto
                edo_futuro = d0;
            end
            
            d11: begin
                cs = 5'b10001;
                rw = 1'b0;
                edo_futuro = d0;
            end
            
            // ... otros estados mantienen l�gica similar
            
            default: begin
                edo_futuro = d0;
                cs = 5'b11110;
            end
        endcase
    end
end

// Proceso 2: Registro de estado - SECUENCIAL
always @(posedge clk or posedge reset) begin
    if (reset) begin
        edo_presente <= d0;
    end else begin
        edo_presente <= edo_futuro;
    end
end

endmodule